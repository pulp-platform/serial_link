// Copyright 2025 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51

`ifndef SERIAL_LINK_REG_SVH
`define SERIAL_LINK_REG_SVH


`define SERIAL_LINK_REG_BASE_ADDR 64'h00000000
`define SERIAL_LINK_REG_SIZE      64'h0000045C


`define SERIAL_LINK_REG_SERIAL_LINK_BASE_ADDR 64'h00000000
`define SERIAL_LINK_REG_SERIAL_LINK_SIZE      64'h0000045C

`define SERIAL_LINK_REG_SERIAL_LINK_CTRL_REG_ADDR   64'h00000000
`define SERIAL_LINK_REG_SERIAL_LINK_CTRL_REG_OFFSET 64'h00000000

`define SERIAL_LINK_REG_SERIAL_LINK_ISOLATED_REG_ADDR   64'h00000004
`define SERIAL_LINK_REG_SERIAL_LINK_ISOLATED_REG_OFFSET 64'h00000004

`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_0_REG_ADDR   64'h00000008
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_0_REG_OFFSET 64'h00000008
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_1_REG_ADDR   64'h0000000C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_1_REG_OFFSET 64'h0000000C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_2_REG_ADDR   64'h00000010
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_2_REG_OFFSET 64'h00000010
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_3_REG_ADDR   64'h00000014
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_3_REG_OFFSET 64'h00000014
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_4_REG_ADDR   64'h00000018
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_4_REG_OFFSET 64'h00000018
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_5_REG_ADDR   64'h0000001C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_5_REG_OFFSET 64'h0000001C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_6_REG_ADDR   64'h00000020
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_6_REG_OFFSET 64'h00000020
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_7_REG_ADDR   64'h00000024
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_7_REG_OFFSET 64'h00000024
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_8_REG_ADDR   64'h00000028
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_8_REG_OFFSET 64'h00000028
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_9_REG_ADDR   64'h0000002C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_9_REG_OFFSET 64'h0000002C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_10_REG_ADDR   64'h00000030
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_10_REG_OFFSET 64'h00000030
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_11_REG_ADDR   64'h00000034
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_11_REG_OFFSET 64'h00000034
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_12_REG_ADDR   64'h00000038
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_12_REG_OFFSET 64'h00000038
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_13_REG_ADDR   64'h0000003C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_13_REG_OFFSET 64'h0000003C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_14_REG_ADDR   64'h00000040
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_14_REG_OFFSET 64'h00000040
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_15_REG_ADDR   64'h00000044
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_15_REG_OFFSET 64'h00000044
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_16_REG_ADDR   64'h00000048
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_16_REG_OFFSET 64'h00000048
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_17_REG_ADDR   64'h0000004C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_17_REG_OFFSET 64'h0000004C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_18_REG_ADDR   64'h00000050
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_18_REG_OFFSET 64'h00000050
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_19_REG_ADDR   64'h00000054
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_19_REG_OFFSET 64'h00000054
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_20_REG_ADDR   64'h00000058
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_20_REG_OFFSET 64'h00000058
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_21_REG_ADDR   64'h0000005C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_21_REG_OFFSET 64'h0000005C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_22_REG_ADDR   64'h00000060
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_22_REG_OFFSET 64'h00000060
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_23_REG_ADDR   64'h00000064
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_23_REG_OFFSET 64'h00000064
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_24_REG_ADDR   64'h00000068
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_24_REG_OFFSET 64'h00000068
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_25_REG_ADDR   64'h0000006C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_25_REG_OFFSET 64'h0000006C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_26_REG_ADDR   64'h00000070
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_26_REG_OFFSET 64'h00000070
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_27_REG_ADDR   64'h00000074
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_27_REG_OFFSET 64'h00000074
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_28_REG_ADDR   64'h00000078
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_28_REG_OFFSET 64'h00000078
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_29_REG_ADDR   64'h0000007C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_29_REG_OFFSET 64'h0000007C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_30_REG_ADDR   64'h00000080
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_30_REG_OFFSET 64'h00000080
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_31_REG_ADDR   64'h00000084
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_31_REG_OFFSET 64'h00000084
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_32_REG_ADDR   64'h00000088
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_32_REG_OFFSET 64'h00000088
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_33_REG_ADDR   64'h0000008C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_33_REG_OFFSET 64'h0000008C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_34_REG_ADDR   64'h00000090
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_34_REG_OFFSET 64'h00000090
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_35_REG_ADDR   64'h00000094
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_35_REG_OFFSET 64'h00000094
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_36_REG_ADDR   64'h00000098
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_36_REG_OFFSET 64'h00000098
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_37_REG_ADDR   64'h0000009C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_DIV_37_REG_OFFSET 64'h0000009C

`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_0_REG_ADDR   64'h000000A0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_0_REG_OFFSET 64'h000000A0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_1_REG_ADDR   64'h000000A4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_1_REG_OFFSET 64'h000000A4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_2_REG_ADDR   64'h000000A8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_2_REG_OFFSET 64'h000000A8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_3_REG_ADDR   64'h000000AC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_3_REG_OFFSET 64'h000000AC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_4_REG_ADDR   64'h000000B0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_4_REG_OFFSET 64'h000000B0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_5_REG_ADDR   64'h000000B4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_5_REG_OFFSET 64'h000000B4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_6_REG_ADDR   64'h000000B8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_6_REG_OFFSET 64'h000000B8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_7_REG_ADDR   64'h000000BC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_7_REG_OFFSET 64'h000000BC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_8_REG_ADDR   64'h000000C0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_8_REG_OFFSET 64'h000000C0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_9_REG_ADDR   64'h000000C4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_9_REG_OFFSET 64'h000000C4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_10_REG_ADDR   64'h000000C8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_10_REG_OFFSET 64'h000000C8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_11_REG_ADDR   64'h000000CC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_11_REG_OFFSET 64'h000000CC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_12_REG_ADDR   64'h000000D0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_12_REG_OFFSET 64'h000000D0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_13_REG_ADDR   64'h000000D4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_13_REG_OFFSET 64'h000000D4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_14_REG_ADDR   64'h000000D8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_14_REG_OFFSET 64'h000000D8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_15_REG_ADDR   64'h000000DC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_15_REG_OFFSET 64'h000000DC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_16_REG_ADDR   64'h000000E0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_16_REG_OFFSET 64'h000000E0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_17_REG_ADDR   64'h000000E4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_17_REG_OFFSET 64'h000000E4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_18_REG_ADDR   64'h000000E8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_18_REG_OFFSET 64'h000000E8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_19_REG_ADDR   64'h000000EC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_19_REG_OFFSET 64'h000000EC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_20_REG_ADDR   64'h000000F0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_20_REG_OFFSET 64'h000000F0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_21_REG_ADDR   64'h000000F4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_21_REG_OFFSET 64'h000000F4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_22_REG_ADDR   64'h000000F8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_22_REG_OFFSET 64'h000000F8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_23_REG_ADDR   64'h000000FC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_23_REG_OFFSET 64'h000000FC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_24_REG_ADDR   64'h00000100
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_24_REG_OFFSET 64'h00000100
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_25_REG_ADDR   64'h00000104
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_25_REG_OFFSET 64'h00000104
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_26_REG_ADDR   64'h00000108
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_26_REG_OFFSET 64'h00000108
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_27_REG_ADDR   64'h0000010C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_27_REG_OFFSET 64'h0000010C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_28_REG_ADDR   64'h00000110
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_28_REG_OFFSET 64'h00000110
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_29_REG_ADDR   64'h00000114
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_29_REG_OFFSET 64'h00000114
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_30_REG_ADDR   64'h00000118
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_30_REG_OFFSET 64'h00000118
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_31_REG_ADDR   64'h0000011C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_31_REG_OFFSET 64'h0000011C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_32_REG_ADDR   64'h00000120
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_32_REG_OFFSET 64'h00000120
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_33_REG_ADDR   64'h00000124
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_33_REG_OFFSET 64'h00000124
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_34_REG_ADDR   64'h00000128
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_34_REG_OFFSET 64'h00000128
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_35_REG_ADDR   64'h0000012C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_35_REG_OFFSET 64'h0000012C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_36_REG_ADDR   64'h00000130
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_36_REG_OFFSET 64'h00000130
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_37_REG_ADDR   64'h00000134
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_START_37_REG_OFFSET 64'h00000134

`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_0_REG_ADDR   64'h00000138
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_0_REG_OFFSET 64'h00000138
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_1_REG_ADDR   64'h0000013C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_1_REG_OFFSET 64'h0000013C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_2_REG_ADDR   64'h00000140
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_2_REG_OFFSET 64'h00000140
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_3_REG_ADDR   64'h00000144
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_3_REG_OFFSET 64'h00000144
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_4_REG_ADDR   64'h00000148
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_4_REG_OFFSET 64'h00000148
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_5_REG_ADDR   64'h0000014C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_5_REG_OFFSET 64'h0000014C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_6_REG_ADDR   64'h00000150
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_6_REG_OFFSET 64'h00000150
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_7_REG_ADDR   64'h00000154
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_7_REG_OFFSET 64'h00000154
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_8_REG_ADDR   64'h00000158
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_8_REG_OFFSET 64'h00000158
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_9_REG_ADDR   64'h0000015C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_9_REG_OFFSET 64'h0000015C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_10_REG_ADDR   64'h00000160
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_10_REG_OFFSET 64'h00000160
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_11_REG_ADDR   64'h00000164
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_11_REG_OFFSET 64'h00000164
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_12_REG_ADDR   64'h00000168
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_12_REG_OFFSET 64'h00000168
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_13_REG_ADDR   64'h0000016C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_13_REG_OFFSET 64'h0000016C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_14_REG_ADDR   64'h00000170
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_14_REG_OFFSET 64'h00000170
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_15_REG_ADDR   64'h00000174
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_15_REG_OFFSET 64'h00000174
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_16_REG_ADDR   64'h00000178
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_16_REG_OFFSET 64'h00000178
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_17_REG_ADDR   64'h0000017C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_17_REG_OFFSET 64'h0000017C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_18_REG_ADDR   64'h00000180
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_18_REG_OFFSET 64'h00000180
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_19_REG_ADDR   64'h00000184
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_19_REG_OFFSET 64'h00000184
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_20_REG_ADDR   64'h00000188
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_20_REG_OFFSET 64'h00000188
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_21_REG_ADDR   64'h0000018C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_21_REG_OFFSET 64'h0000018C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_22_REG_ADDR   64'h00000190
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_22_REG_OFFSET 64'h00000190
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_23_REG_ADDR   64'h00000194
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_23_REG_OFFSET 64'h00000194
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_24_REG_ADDR   64'h00000198
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_24_REG_OFFSET 64'h00000198
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_25_REG_ADDR   64'h0000019C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_25_REG_OFFSET 64'h0000019C
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_26_REG_ADDR   64'h000001A0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_26_REG_OFFSET 64'h000001A0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_27_REG_ADDR   64'h000001A4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_27_REG_OFFSET 64'h000001A4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_28_REG_ADDR   64'h000001A8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_28_REG_OFFSET 64'h000001A8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_29_REG_ADDR   64'h000001AC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_29_REG_OFFSET 64'h000001AC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_30_REG_ADDR   64'h000001B0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_30_REG_OFFSET 64'h000001B0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_31_REG_ADDR   64'h000001B4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_31_REG_OFFSET 64'h000001B4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_32_REG_ADDR   64'h000001B8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_32_REG_OFFSET 64'h000001B8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_33_REG_ADDR   64'h000001BC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_33_REG_OFFSET 64'h000001BC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_34_REG_ADDR   64'h000001C0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_34_REG_OFFSET 64'h000001C0
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_35_REG_ADDR   64'h000001C4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_35_REG_OFFSET 64'h000001C4
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_36_REG_ADDR   64'h000001C8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_36_REG_OFFSET 64'h000001C8
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_37_REG_ADDR   64'h000001CC
`define SERIAL_LINK_REG_SERIAL_LINK_TX_PHY_CLK_END_37_REG_OFFSET 64'h000001CC

`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_EN_REG_ADDR   64'h000001D0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_EN_REG_OFFSET 64'h000001D0

`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_CH_SEL_REG_ADDR   64'h000001D4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_CH_SEL_REG_OFFSET 64'h000001D4

`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_0_REG_ADDR   64'h000001D8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_0_REG_OFFSET 64'h000001D8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_1_REG_ADDR   64'h000001DC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_1_REG_OFFSET 64'h000001DC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_2_REG_ADDR   64'h000001E0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_2_REG_OFFSET 64'h000001E0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_3_REG_ADDR   64'h000001E4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_3_REG_OFFSET 64'h000001E4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_4_REG_ADDR   64'h000001E8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_4_REG_OFFSET 64'h000001E8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_5_REG_ADDR   64'h000001EC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_5_REG_OFFSET 64'h000001EC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_6_REG_ADDR   64'h000001F0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_6_REG_OFFSET 64'h000001F0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_7_REG_ADDR   64'h000001F4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_7_REG_OFFSET 64'h000001F4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_8_REG_ADDR   64'h000001F8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_8_REG_OFFSET 64'h000001F8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_9_REG_ADDR   64'h000001FC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_9_REG_OFFSET 64'h000001FC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_10_REG_ADDR   64'h00000200
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_10_REG_OFFSET 64'h00000200
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_11_REG_ADDR   64'h00000204
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_11_REG_OFFSET 64'h00000204
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_12_REG_ADDR   64'h00000208
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_12_REG_OFFSET 64'h00000208
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_13_REG_ADDR   64'h0000020C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_13_REG_OFFSET 64'h0000020C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_14_REG_ADDR   64'h00000210
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_14_REG_OFFSET 64'h00000210
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_15_REG_ADDR   64'h00000214
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_15_REG_OFFSET 64'h00000214
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_16_REG_ADDR   64'h00000218
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_16_REG_OFFSET 64'h00000218
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_17_REG_ADDR   64'h0000021C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_17_REG_OFFSET 64'h0000021C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_18_REG_ADDR   64'h00000220
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_18_REG_OFFSET 64'h00000220
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_19_REG_ADDR   64'h00000224
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_19_REG_OFFSET 64'h00000224
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_20_REG_ADDR   64'h00000228
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_20_REG_OFFSET 64'h00000228
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_21_REG_ADDR   64'h0000022C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_21_REG_OFFSET 64'h0000022C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_22_REG_ADDR   64'h00000230
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_22_REG_OFFSET 64'h00000230
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_23_REG_ADDR   64'h00000234
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_23_REG_OFFSET 64'h00000234
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_24_REG_ADDR   64'h00000238
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_24_REG_OFFSET 64'h00000238
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_25_REG_ADDR   64'h0000023C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_25_REG_OFFSET 64'h0000023C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_26_REG_ADDR   64'h00000240
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_26_REG_OFFSET 64'h00000240
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_27_REG_ADDR   64'h00000244
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_27_REG_OFFSET 64'h00000244
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_28_REG_ADDR   64'h00000248
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_28_REG_OFFSET 64'h00000248
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_29_REG_ADDR   64'h0000024C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_29_REG_OFFSET 64'h0000024C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_30_REG_ADDR   64'h00000250
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_30_REG_OFFSET 64'h00000250
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_31_REG_ADDR   64'h00000254
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_31_REG_OFFSET 64'h00000254
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_32_REG_ADDR   64'h00000258
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_32_REG_OFFSET 64'h00000258
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_33_REG_ADDR   64'h0000025C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_33_REG_OFFSET 64'h0000025C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_34_REG_ADDR   64'h00000260
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_34_REG_OFFSET 64'h00000260
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_35_REG_ADDR   64'h00000264
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_35_REG_OFFSET 64'h00000264
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_36_REG_ADDR   64'h00000268
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_36_REG_OFFSET 64'h00000268
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_37_REG_ADDR   64'h0000026C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_37_REG_OFFSET 64'h0000026C

`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_REG_ADDR   64'h00000270
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_IN_DATA_REG_OFFSET 64'h00000270

`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_0_REG_ADDR   64'h00000274
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_0_REG_OFFSET 64'h00000274
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_1_REG_ADDR   64'h00000278
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_1_REG_OFFSET 64'h00000278
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_2_REG_ADDR   64'h0000027C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_2_REG_OFFSET 64'h0000027C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_3_REG_ADDR   64'h00000280
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_3_REG_OFFSET 64'h00000280
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_4_REG_ADDR   64'h00000284
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_4_REG_OFFSET 64'h00000284
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_5_REG_ADDR   64'h00000288
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_5_REG_OFFSET 64'h00000288
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_6_REG_ADDR   64'h0000028C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_6_REG_OFFSET 64'h0000028C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_7_REG_ADDR   64'h00000290
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_7_REG_OFFSET 64'h00000290
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_8_REG_ADDR   64'h00000294
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_8_REG_OFFSET 64'h00000294
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_9_REG_ADDR   64'h00000298
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_9_REG_OFFSET 64'h00000298
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_10_REG_ADDR   64'h0000029C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_10_REG_OFFSET 64'h0000029C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_11_REG_ADDR   64'h000002A0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_11_REG_OFFSET 64'h000002A0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_12_REG_ADDR   64'h000002A4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_12_REG_OFFSET 64'h000002A4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_13_REG_ADDR   64'h000002A8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_13_REG_OFFSET 64'h000002A8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_14_REG_ADDR   64'h000002AC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_14_REG_OFFSET 64'h000002AC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_15_REG_ADDR   64'h000002B0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_15_REG_OFFSET 64'h000002B0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_16_REG_ADDR   64'h000002B4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_16_REG_OFFSET 64'h000002B4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_17_REG_ADDR   64'h000002B8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_17_REG_OFFSET 64'h000002B8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_18_REG_ADDR   64'h000002BC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_18_REG_OFFSET 64'h000002BC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_19_REG_ADDR   64'h000002C0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_19_REG_OFFSET 64'h000002C0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_20_REG_ADDR   64'h000002C4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_20_REG_OFFSET 64'h000002C4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_21_REG_ADDR   64'h000002C8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_21_REG_OFFSET 64'h000002C8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_22_REG_ADDR   64'h000002CC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_22_REG_OFFSET 64'h000002CC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_23_REG_ADDR   64'h000002D0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_23_REG_OFFSET 64'h000002D0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_24_REG_ADDR   64'h000002D4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_24_REG_OFFSET 64'h000002D4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_25_REG_ADDR   64'h000002D8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_25_REG_OFFSET 64'h000002D8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_26_REG_ADDR   64'h000002DC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_26_REG_OFFSET 64'h000002DC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_27_REG_ADDR   64'h000002E0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_27_REG_OFFSET 64'h000002E0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_28_REG_ADDR   64'h000002E4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_28_REG_OFFSET 64'h000002E4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_29_REG_ADDR   64'h000002E8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_29_REG_OFFSET 64'h000002E8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_30_REG_ADDR   64'h000002EC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_30_REG_OFFSET 64'h000002EC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_31_REG_ADDR   64'h000002F0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_31_REG_OFFSET 64'h000002F0
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_32_REG_ADDR   64'h000002F4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_32_REG_OFFSET 64'h000002F4
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_33_REG_ADDR   64'h000002F8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_33_REG_OFFSET 64'h000002F8
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_34_REG_ADDR   64'h000002FC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_34_REG_OFFSET 64'h000002FC
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_35_REG_ADDR   64'h00000300
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_35_REG_OFFSET 64'h00000300
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_36_REG_ADDR   64'h00000304
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_36_REG_OFFSET 64'h00000304
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_37_REG_ADDR   64'h00000308
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_37_REG_OFFSET 64'h00000308

`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_REG_ADDR   64'h0000030C
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_REG_OFFSET 64'h0000030C

`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_CTRL_REG_ADDR   64'h00000310
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_CTRL_REG_OFFSET 64'h00000310

`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_EN_REG_ADDR   64'h00000314
`define SERIAL_LINK_REG_SERIAL_LINK_RAW_MODE_OUT_EN_REG_OFFSET 64'h00000314

`define SERIAL_LINK_REG_SERIAL_LINK_FLOW_CONTROL_FIFO_CLEAR_REG_ADDR   64'h00000318
`define SERIAL_LINK_REG_SERIAL_LINK_FLOW_CONTROL_FIFO_CLEAR_REG_OFFSET 64'h00000318

`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CFG_REG_ADDR   64'h0000031C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CFG_REG_OFFSET 64'h0000031C

`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_0_REG_ADDR   64'h00000320
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_0_REG_OFFSET 64'h00000320
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_1_REG_ADDR   64'h00000324
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_1_REG_OFFSET 64'h00000324
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_2_REG_ADDR   64'h00000328
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_2_REG_OFFSET 64'h00000328
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_3_REG_ADDR   64'h0000032C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_3_REG_OFFSET 64'h0000032C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_4_REG_ADDR   64'h00000330
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_4_REG_OFFSET 64'h00000330
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_5_REG_ADDR   64'h00000334
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_5_REG_OFFSET 64'h00000334
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_6_REG_ADDR   64'h00000338
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_6_REG_OFFSET 64'h00000338
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_7_REG_ADDR   64'h0000033C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_7_REG_OFFSET 64'h0000033C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_8_REG_ADDR   64'h00000340
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_8_REG_OFFSET 64'h00000340
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_9_REG_ADDR   64'h00000344
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_9_REG_OFFSET 64'h00000344
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_10_REG_ADDR   64'h00000348
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_10_REG_OFFSET 64'h00000348
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_11_REG_ADDR   64'h0000034C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_11_REG_OFFSET 64'h0000034C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_12_REG_ADDR   64'h00000350
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_12_REG_OFFSET 64'h00000350
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_13_REG_ADDR   64'h00000354
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_13_REG_OFFSET 64'h00000354
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_14_REG_ADDR   64'h00000358
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_14_REG_OFFSET 64'h00000358
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_15_REG_ADDR   64'h0000035C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_15_REG_OFFSET 64'h0000035C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_16_REG_ADDR   64'h00000360
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_16_REG_OFFSET 64'h00000360
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_17_REG_ADDR   64'h00000364
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_17_REG_OFFSET 64'h00000364
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_18_REG_ADDR   64'h00000368
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_18_REG_OFFSET 64'h00000368
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_19_REG_ADDR   64'h0000036C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_19_REG_OFFSET 64'h0000036C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_20_REG_ADDR   64'h00000370
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_20_REG_OFFSET 64'h00000370
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_21_REG_ADDR   64'h00000374
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_21_REG_OFFSET 64'h00000374
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_22_REG_ADDR   64'h00000378
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_22_REG_OFFSET 64'h00000378
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_23_REG_ADDR   64'h0000037C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_23_REG_OFFSET 64'h0000037C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_24_REG_ADDR   64'h00000380
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_24_REG_OFFSET 64'h00000380
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_25_REG_ADDR   64'h00000384
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_25_REG_OFFSET 64'h00000384
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_26_REG_ADDR   64'h00000388
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_26_REG_OFFSET 64'h00000388
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_27_REG_ADDR   64'h0000038C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_27_REG_OFFSET 64'h0000038C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_28_REG_ADDR   64'h00000390
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_28_REG_OFFSET 64'h00000390
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_29_REG_ADDR   64'h00000394
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_29_REG_OFFSET 64'h00000394
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_30_REG_ADDR   64'h00000398
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_30_REG_OFFSET 64'h00000398
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_31_REG_ADDR   64'h0000039C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_31_REG_OFFSET 64'h0000039C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_32_REG_ADDR   64'h000003A0
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_32_REG_OFFSET 64'h000003A0
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_33_REG_ADDR   64'h000003A4
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_33_REG_OFFSET 64'h000003A4
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_34_REG_ADDR   64'h000003A8
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_34_REG_OFFSET 64'h000003A8
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_35_REG_ADDR   64'h000003AC
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_35_REG_OFFSET 64'h000003AC
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_36_REG_ADDR   64'h000003B0
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_36_REG_OFFSET 64'h000003B0
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_37_REG_ADDR   64'h000003B4
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_37_REG_OFFSET 64'h000003B4

`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CTRL_REG_ADDR   64'h000003B8
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CTRL_REG_OFFSET 64'h000003B8

`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CFG_REG_ADDR   64'h000003BC
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CFG_REG_OFFSET 64'h000003BC

`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CTRL_REG_ADDR   64'h000003C0
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CTRL_REG_OFFSET 64'h000003C0

`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_0_REG_ADDR   64'h000003C4
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_0_REG_OFFSET 64'h000003C4
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_1_REG_ADDR   64'h000003C8
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_1_REG_OFFSET 64'h000003C8
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_2_REG_ADDR   64'h000003CC
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_2_REG_OFFSET 64'h000003CC
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_3_REG_ADDR   64'h000003D0
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_3_REG_OFFSET 64'h000003D0
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_4_REG_ADDR   64'h000003D4
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_4_REG_OFFSET 64'h000003D4
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_5_REG_ADDR   64'h000003D8
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_5_REG_OFFSET 64'h000003D8
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_6_REG_ADDR   64'h000003DC
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_6_REG_OFFSET 64'h000003DC
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_7_REG_ADDR   64'h000003E0
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_7_REG_OFFSET 64'h000003E0
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_8_REG_ADDR   64'h000003E4
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_8_REG_OFFSET 64'h000003E4
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_9_REG_ADDR   64'h000003E8
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_9_REG_OFFSET 64'h000003E8
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_10_REG_ADDR   64'h000003EC
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_10_REG_OFFSET 64'h000003EC
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_11_REG_ADDR   64'h000003F0
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_11_REG_OFFSET 64'h000003F0
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_12_REG_ADDR   64'h000003F4
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_12_REG_OFFSET 64'h000003F4
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_13_REG_ADDR   64'h000003F8
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_13_REG_OFFSET 64'h000003F8
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_14_REG_ADDR   64'h000003FC
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_14_REG_OFFSET 64'h000003FC
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_15_REG_ADDR   64'h00000400
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_15_REG_OFFSET 64'h00000400
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_16_REG_ADDR   64'h00000404
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_16_REG_OFFSET 64'h00000404
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_17_REG_ADDR   64'h00000408
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_17_REG_OFFSET 64'h00000408
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_18_REG_ADDR   64'h0000040C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_18_REG_OFFSET 64'h0000040C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_19_REG_ADDR   64'h00000410
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_19_REG_OFFSET 64'h00000410
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_20_REG_ADDR   64'h00000414
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_20_REG_OFFSET 64'h00000414
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_21_REG_ADDR   64'h00000418
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_21_REG_OFFSET 64'h00000418
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_22_REG_ADDR   64'h0000041C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_22_REG_OFFSET 64'h0000041C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_23_REG_ADDR   64'h00000420
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_23_REG_OFFSET 64'h00000420
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_24_REG_ADDR   64'h00000424
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_24_REG_OFFSET 64'h00000424
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_25_REG_ADDR   64'h00000428
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_25_REG_OFFSET 64'h00000428
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_26_REG_ADDR   64'h0000042C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_26_REG_OFFSET 64'h0000042C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_27_REG_ADDR   64'h00000430
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_27_REG_OFFSET 64'h00000430
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_28_REG_ADDR   64'h00000434
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_28_REG_OFFSET 64'h00000434
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_29_REG_ADDR   64'h00000438
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_29_REG_OFFSET 64'h00000438
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_30_REG_ADDR   64'h0000043C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_30_REG_OFFSET 64'h0000043C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_31_REG_ADDR   64'h00000440
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_31_REG_OFFSET 64'h00000440
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_32_REG_ADDR   64'h00000444
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_32_REG_OFFSET 64'h00000444
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_33_REG_ADDR   64'h00000448
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_33_REG_OFFSET 64'h00000448
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_34_REG_ADDR   64'h0000044C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_34_REG_OFFSET 64'h0000044C
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_35_REG_ADDR   64'h00000450
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_35_REG_OFFSET 64'h00000450
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_36_REG_ADDR   64'h00000454
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_36_REG_OFFSET 64'h00000454
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_37_REG_ADDR   64'h00000458
`define SERIAL_LINK_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_37_REG_OFFSET 64'h00000458


`endif /* SERIAL_LINK_REG_SVH */
