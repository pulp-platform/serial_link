`ifndef SERIAL_LINK_SINGLE_CHANNEL_REG_SVH
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SVH


`define SERIAL_LINK_SINGLE_CHANNEL_REG_BASE_ADDR 64'h00000000
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SIZE      64'h00000050


`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_BASE_ADDR 64'h00000000
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_SIZE      64'h00000050

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CTRL_REG_ADDR   64'h00000000
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CTRL_REG_OFFSET 64'h00000000

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_ISOLATED_REG_ADDR   64'h00000004
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_ISOLATED_REG_OFFSET 64'h00000004

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_DIV_0_REG_ADDR   64'h00000008
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_DIV_0_REG_OFFSET 64'h00000008

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_START_0_REG_ADDR   64'h0000000C
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_START_0_REG_OFFSET 64'h0000000C

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_END_0_REG_ADDR   64'h00000010
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_END_0_REG_OFFSET 64'h00000010

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_EN_REG_ADDR   64'h00000014
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_EN_REG_OFFSET 64'h00000014

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_CH_SEL_REG_ADDR   64'h00000018
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_CH_SEL_REG_OFFSET 64'h00000018

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_0_REG_ADDR   64'h0000001C
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_0_REG_OFFSET 64'h0000001C

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_DATA_REG_ADDR   64'h00000020
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_DATA_REG_OFFSET 64'h00000020

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_0_REG_ADDR   64'h00000024
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_0_REG_OFFSET 64'h00000024

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_REG_ADDR   64'h00000028
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_REG_OFFSET 64'h00000028

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_CTRL_REG_ADDR   64'h0000002C
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_CTRL_REG_OFFSET 64'h0000002C

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_EN_REG_ADDR   64'h00000030
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_EN_REG_OFFSET 64'h00000030

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_FLOW_CONTROL_FIFO_CLEAR_REG_ADDR   64'h00000034
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_FLOW_CONTROL_FIFO_CLEAR_REG_OFFSET 64'h00000034

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CFG_REG_ADDR   64'h00000038
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CFG_REG_OFFSET 64'h00000038

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_0_REG_ADDR   64'h0000003C
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CH_EN_0_REG_OFFSET 64'h0000003C

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CTRL_REG_ADDR   64'h00000040
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_TX_CTRL_REG_OFFSET 64'h00000040

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CFG_REG_ADDR   64'h00000044
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CFG_REG_OFFSET 64'h00000044

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CTRL_REG_ADDR   64'h00000048
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CTRL_REG_OFFSET 64'h00000048

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_0_REG_ADDR   64'h0000004C
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CHANNEL_ALLOC_RX_CH_EN_0_REG_OFFSET 64'h0000004C


`endif /* SERIAL_LINK_SINGLE_CHANNEL_REG_SVH */
