// Copyright 2025 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51

`ifndef SERIAL_LINK_SINGLE_CHANNEL_REG_SVH
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SVH


`define SERIAL_LINK_SINGLE_CHANNEL_REG_BASE_ADDR 64'h00000000
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SIZE      64'h00000804


`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_BASE_ADDR 64'h00000000
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_SIZE      64'h00000804

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CTRL_REG_ADDR   64'h00000000
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_CTRL_REG_OFFSET 64'h00000000

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_ISOLATED_REG_ADDR   64'h00000004
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_ISOLATED_REG_OFFSET 64'h00000004

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_EN_REG_ADDR   64'h00000008
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_EN_REG_OFFSET 64'h00000008

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_DATA_REG_ADDR   64'h0000000C
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_DATA_REG_OFFSET 64'h0000000C

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_CH_SEL_REG_ADDR   64'h00000010
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_CH_SEL_REG_OFFSET 64'h00000010

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_REG_ADDR   64'h00000014
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_REG_OFFSET 64'h00000014

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_CTRL_REG_ADDR   64'h00000018
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_DATA_FIFO_CTRL_REG_OFFSET 64'h00000018

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_EN_REG_ADDR   64'h0000001C
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_EN_REG_OFFSET 64'h0000001C

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_FLOW_CONTROL_FIFO_CLEAR_REG_ADDR   64'h00000020
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_FLOW_CONTROL_FIFO_CLEAR_REG_OFFSET 64'h00000020

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_0_REG_ADDR   64'h00000100
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_IN_DATA_VALID_0_REG_OFFSET 64'h00000100

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_0_REG_ADDR   64'h00000200
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_RAW_MODE_OUT_CH_MASK_0_REG_OFFSET 64'h00000200

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_DIV_0_REG_ADDR   64'h00000300
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_DIV_0_REG_OFFSET 64'h00000300

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_START_0_REG_ADDR   64'h00000400
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_START_0_REG_OFFSET 64'h00000400

`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_END_0_REG_ADDR   64'h00000500
`define SERIAL_LINK_SINGLE_CHANNEL_REG_SERIAL_LINK_TX_PHY_CLK_END_0_REG_OFFSET 64'h00000500


`endif /* SERIAL_LINK_SINGLE_CHANNEL_REG_SVH */
